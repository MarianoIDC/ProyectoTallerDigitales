module ROM_Ins
#(
    parameter 
                 addr_bits = 8, // required bits to store 16 elements
                 data_width = 32 // each element has 1-bit Background or Image
)
(
    input logic [addr_bits-1:0] addr,
    output reg [data_width-1:0] data  
);
always @*
	begin
		 case(addr)
				8'b00000000 : data = 32'he3a00b01;//0 Guardar en memoria la frase
				8'b00000001 : data = 32'he3a01c05;//1 Guardar los datos descifrados
				8'b00000010 : data = 32'he3a0b002;//2 escoger desencriptado
				8'b00000011 : data = 32'he3a0207d;//3 m
				8'b00000100 : data = 32'he4802004;//4 s
				8'b00000101 : data = 32'he3a02050;//5 m
				8'b00000110 : data = 32'he4802004;//6 s
				8'b00000111 : data = 32'he3a02059;//7 m
				8'b00001000 : data = 32'he4802004;//8 s 
				8'b00001001 : data = 32'he3a02059;//9
				8'b00001010 : data = 32'he4802004;//10
				8'b00001011 : data = 32'he3a0205a;//11
				8'b00001100 : data = 32'he4802004;//12
				8'b00001101 : data = 32'he3a02019;//13
				8'b00001110 : data = 32'he4802004;//14 ///////////
				8'b00001111 : data = 32'he3a02015;//15
				8'b00010000 : data = 32'he4802004;//16
				8'b00010001 : data = 32'he3a02062;//17
				8'b00010010 : data = 32'he4802004;//18
				8'b00010011 : data = 32'he3a0205a;//19
				8'b00010100 : data = 32'he4802004;//20
				8'b00010101 : data = 32'he3a02047;//21
				8'b00010110 : data = 32'he4802004;//22
				8'b00010111 : data = 32'he3a02059;//23
				8'b00011000 : data = 32'he4802004;//24
				8'b00011001 : data = 32'he3a02051;//25
				8'b00011010 : data = 32'he4802004;//26
				8'b00011011 : data = 32'he3a02014;//27
				8'b00011100 : data = 32'he4802004;//28
				8'b00011101 : data = 32'he3a0200a;//29
				8'b00011110 : data = 32'he4802004;//30////////////////
				8'b00011111 : data = 32'he3a00b01;//31  Esta bien
				8'b00100000 : data = 32'he1a02000;//32
				8'b00100001 : data = 32'he1a07001;//33
				8'b00100010 : data = 32'he35b0001;//34
				8'b00100011 : data = 32'h0a000003;//35
				8'b00100100 : data = 32'he35b0002;//36
				8'b00100101 : data = 32'h0a00000b;//37
				8'b00100110 : data = 32'he35b0003;//38
				8'b00100111 : data = 32'h0a000013;//39
				8'b00101000 : data = 32'he4903004;//40
				8'b00101001 : data = 32'he353000a;//41
				8'b00101010 : data = 32'h1a000000;//42
				8'b00101011 : data = 32'hea000018;//43
				8'b00101100 : data = 32'he3a09035;//44
				8'b00101101 : data = 32'he4914004;//45
				8'b00101110 : data = 32'he4925004;//46
				8'b00101111 : data = 32'he0296005;//47
				8'b00110000 : data = 32'he4876004;//48
				8'b00110001 : data = 32'heafffff5;//49
				8'b00110010 : data = 32'he4903004;//50
				8'b00110011 : data = 32'he353000a;//51
				8'b00110100 : data = 32'h1a000000;//52
				8'b00110101 : data = 32'hea00000e;//53
				8'b00110110 : data = 32'he3a090ff;//54
				8'b00110111 : data = 32'he4914004;//55
				8'b00111000 : data = 32'he4925004;//56
				8'b00111001 : data = 32'he0496005;//57
				8'b00111010 : data = 32'he4876004;//58
				8'b00111011 : data = 32'heafffff5;//59
				8'b00111100 : data = 32'he4903004;//60
				8'b00111101 : data = 32'he353000a;//61
				8'b00111110 : data = 32'h1a000000;//62
				8'b00111111 : data = 32'hea000004;//63
				8'b01000000 : data = 32'he4914004;//64
				8'b01000001 : data = 32'he4925004;//65
				8'b01000010 : data = 32'he2856002;//66
				8'b01000011 : data = 32'he4876004;//67
				8'b01000100 : data = 32'heafffff6;//68
				8'b01000101 : data = 32'h00000000;//69
		
			  default   : data = 32'b00000000000000000000000000000000; // 15
		 endcase 
	end
endmodule 